interface adder_if(input logic clk, reset);
  logic [3:0] a;
  logic [3:0] b;
  logic [4:0] y;
endinterface
/*
interface add_if(input logic clk, reset);
  logic [7:0] ip1, ip2;
  logic [8:0] out;
endinterface*/
  
