package adder_pkg;
   import uvm_pkg::*;
   `include "uvm_macros.svh"
   //`include "simpleadder_configuration.svh"
   `include "seq_item.sv"
   `include "sequence.sv"
   `include "driver.sv" 
   `include "monitor.sv"
   `include "agent.sv"
  // `include "simpleadder_scoreboard.svh"
   `include "env.sv"
   `include "test.sv"
endpackage
